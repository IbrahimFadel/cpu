`define READ 0
`define WRITE 1

`define NO_RESET 0
`define YES_RESET 1

`define READ_SEL_PC 0
`define READ_SEL_DB 1
`define READ_SEL_AR 2

`define AR_READ_PC 0
`define AR_READ_DST_REG 1

`define INT_DATA_READ_PC 0
`define INT_DATA_READ_REG 1