`define R0 8'h0
`define R1 8'h1
`define R2 8'h2
`define R3 8'h3
