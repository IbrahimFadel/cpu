`define MOV_REG_REG 8'h0
`define MOV_REG_LIT 8'h1
`define MOV_REG_MEM 8'h2
`define MOV_MEM_REG 8'h3

`define ADD_REG_LIT 8'h4

`define OP_ADD 4'h0

`define R0 8'h0
`define R1 8'h1
`define R2 8'h2
`define R3 8'h3

`define RESET 1'b0
`define NO_RESET 1'b1
