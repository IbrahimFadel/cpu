parameter WORD_SIZE = 32,
parameter NUM_REG = 32,
parameter ADDRESS_SIZE = 9
