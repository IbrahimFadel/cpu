module alu ();

endmodule
