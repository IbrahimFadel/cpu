`define FETCH1 1
`define FETCH2 2

`define MOV_REG_REG1 3