`define BYTE_SIZE 8
`define WORD_SIZE 16
`define ROM_SIZE 256
`define RAM_SIZE 256
